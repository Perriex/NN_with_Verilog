`timescale 1ns/1ns

module Controller();

    parameter size = 16;

endmodule